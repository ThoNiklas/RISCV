//`define TB
