module RISCV #(parameter REG_BITS=32, parameter ADDR_BITS=5) 
(
    input logic CLK, RST
);

    ProgramCounter #(.REG_BITS(REG_BITS)) programCounter (.clk(c 

endmodule

