module ExtendImm #(parameter REG_BITS=32)
(
    input logic [24:0] in,
    output logic [REG_BITS-1:0] out
);

endmodule

