module ExtendResult #(parameter REG_BITS=32)
(
    input logic [REG_BITS-1:0] in,
    output logic [REG_BITS-1:0] out
);

endmodule

