//`define TESTBENCH 
