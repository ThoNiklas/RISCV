`define TESTBENCH
